{"table_done": ["ATT_MID_CHA_TRAN_PD_TEMP", "CONSUMERACTUALMAP", "CSTCONSUMERACTUALBET_V", "DATABLOCK", "DATAMODLE", "DATA_ID_MAP_INFO", "DX_WMY", "ISC_PMS_DEPT", "ISC_PMS_IS_USER", "ISC_SPECIALORG_UNIT_LOCEXT", "ISC_SPECIALORG_UNIT_LOCEXT0802", "ISC_SYSCHRO_LOG", "ISC_USER_LOCEXT", "ISC_USER_LOCEXT0802SF", "MV_ZH_BZQX_QUERY", "MV_ZH_PWBZQX_QUERY", "OBJECTPOOL", "OPC_CODE", "OPC_CONFINFO", "OPC_MANAGER", "OPC_MODEL", "OPC_MODEL_COLS", "OPC_MODEL_COLS20151218", "PMS_JB_GXJL", "SERVERCONFIG", "SERVERMANAGERCONFIG", "TEST", "T_CMS_C_METER_MP_RELA", "T_CMS_C_MP", "T_CMS_G_KK", "T_CMS_G_TRAN", "T_CMS_G_TRAN0422", "T_CMS_G_TRAN0810", "T_CMS_G_TRAN1009", "T_CMS_G_TRAN2016034", "T_CMS_G_TRAN_BAK", "T_CMS_G_TRAN_CLH", "T_CMS_IT_RUM", "T_CMS_METER_MP_RELA", "T_CMS_MP_IT_RELA", "T_CMS_R_COLL_OBJ", "T_CMS_USERDOC_CHECK_LIST", "T_DTOOLS_DRRZ", "T_DTOOLS_IMPEXP_LX", "T_DTOOLS_IMPEXP_ZDPZ", "T_DW_BZZX_BHGNFL", "T_DW_BZZX_BZBGSQD", "T_DW_BZZX_BZFLB", "T_DW_BZZX_BZSJBGHZ", "T_DW_BZZX_BZSJBGHZ_BAK", "T_DW_BZZX_BZSJBGJL", "T_DW_BZZX_BZSJBGJL_BAK", "T_DW_BZZX_CJSBLX", "T_DW_BZZX_GGDMB", "T_DW_BZZX_GNWZBM", "T_DW_BZZX_GZQXYYDM", "T_DW_BZZX_ORDER", "T_DW_BZZX_SBBZCSMB", "T_DW_BZZX_SBFL", "T_DW_BZZX_SBXHB", "T_DW_BZZX_SBXHBZCSB", "T_DW_BZZX_SBXHBZCSB_VER", "T_DW_BZZX_SBXHB_BAK", "T_DW_BZZX_SBXHB_BF", "T_DW_BZZX_SBXHB_BFB", "T_DW_BZZX_SBXHB_VER", "T_DW_BZZX_SBXHB_ZJ_TEMP", "T_DW_BZZX_SCCJ", "T_DW_BZZX_SCCJ_BDSJ_BF", "T_DW_BZZX_SCCJ_BDSJ_DEL", "T_DW_BZZX_SCCJ_BF", "T_DW_BZZX_SCCJ_GFSJ_TEMP", "T_DW_BZZX_SCCJ_HBSJ_TEMP", "T_DW_BZZX_SCCJ_VER", "T_DW_CIMSVG_CITY_CFG", "T_DW_CIMSVG_CONFIG", "T_DW_DDZZJG", "T_DW_DWZY_PWGM", "T_DW_FZBBB_BDRL", "T_DW_FZBBB_JLXL", "T_DW_JK_ERPSERVICENAME", "T_DW_JK_GNWZ", "T_DW_JK_IMS_CONFIG", "T_DW_JK_IMS_DEPART", "T_DW_JK_IMS_JKZBINFO", "T_DW_JK_JHBPZ", "T_DW_JK_JHBSXPZ", "T_DW_JK_JLDGX", "T_DW_JK_YKBZ_TXSH", "T_DW_PZ_TYXH_FW_TEMP", "T_DW_QJ_CBDE", "T_DW_QJ_CFDD", "T_DW_QJ_SYGHJL", "T_DW_QJ_ZTB", "T_DW_SBBG_BGSBLB", "T_DW_SBBG_BGSBQD", "CSTEUQCONSUMER_V", "T_DW_SBBG_DMSMESSAGELOG", "T_DW_SBBG_GCBHPZ", "T_DW_SBBG_RWGL", "T_DW_SBBG_SBBGSQD_SHXX", "T_DW_SBBG_SBBGSQD", "over_view", "T_ZH_BDJYH_PJXMJG", "T_DW_ZCGL_SWZCBB_BFCY_2", "T_SB_PZ_JMXX", "T_ZH_YJJX_ZBZSDWPZ", "T_ZH_JGDY_JGXJXMZB", "T_TD_EXT_LOG_JOBOPERATION", "T_YJ_ZXGL_OMSDLXX", "T_ZH_YJJX_KHDWPZ", "T_YJ_DWYJ_BZHZY_ZYWB_GGYS", "T_YJ_GGSJ_DMFL", "T_YJ_DWYJ_ERPSERVICE", "T_ZH_ZTJX_PDPJRWBGGL", "T_EDC_BUFF_GL", "T_ZH_JSJD_JDHDXZGL", "T_ZH_GYSPJ_GZXX", "T_ZH_JGGL_JGXMJYZB", "T_TD_EXT_JOB_ANALYSIS", "T_ZH_JSJD_PJXZ", "T_ZH_YJJX_JSXZXJG", "T_SB_ZNYC_DLQ", "T_ZH_JGGL_JGXMBZB", "T_MXPMS_WEBSERVICE_ROUTE", "T_MXPMS_WORKITEM_READ", "T_SB_ZNYC_KZCS_DY", "T_ZH_BDJYH_PJSB", "T_ZH_BDDDJC_JCJH", "T_ZH_ZTJX_XLDYKFQZB", "T_PWGC_ZRC", "T_ZHJH_JGDX_XXJDZB", "T_SB_ZWYC_DLZD", "T_YJ_DWYJ_BZHZY_ZYWB_XSNR", "T_SB_ZWYC_ZSDRQ_VER", "T_SB_ZNYC_DLDRQ", "T_YJ_FC_CONS_CERT_RELA", "T_PWGC_PWZXGCGL_ZXDX_TZ_TMP", "T_PWGC_XMCBK_DBXM_DR", "T_XB_PWYW_PMS_ZTJC", "T_YJ_DWYJ_BZHZY_ZYWB_SYML", "T_YJ_GZQX_GDZPTREE", "T_PWGC_WZFWGYS", "T_SB_ZNYC_PDBYQ", "T_ZH_ZTJX_BDPJRW", "T_YJ_DWYJ_DDZY_PWDLBTDZYQKTJB", "T_ZH_JSJD_JSJDBZ", "T_PWGC_PWXQ_FXTZZB_TMP", "T_ZH_ZTJX_ZTLXXD", "T_ZH_JGDX_IN_TAB", "T_SB_SCFZSS_ZMXT", "T_PWGC_PWXQ_GJCXZB", "T_YJ_DWYJ_BZSYM_RYJSB", "T_SB_PZ_PMSERPTABLE", "T_YJ_JCZX_ZHBBGL_DLSBFJHTYBB", "T_ZH_DXGL_XXJDGZGMTJB", "T_SB_ZWYC_DKX_VER", "T_PWGC_FYXMHZTJ", "T_MXPMS_WORKFLOW_LOG", "over_view"], "pms": [""]}